`timescale 1ns/1ns
`include "orgatefinal.v"
module orgatefinal_tb;
reg [3:0]in;
wire f;
orgatefinal ogf(in,f);
initial
begin
$dumpfile("orgatefinal_tb.vcd");
$dumpvars(0,orgatefinal_tb);

        in = 4'b0000; #20;
        in = 4'b0001; #20;
        in = 4'b0010; #20;
        in = 4'b0011; #20;
        in = 4'b0100; #20;
        in = 4'b0101; #20;
        in = 4'b0110; #20;
        in = 4'b0111; #20;
        in = 4'b1000; #20;
        in = 4'b1001; #20;
        in = 4'b1010; #20;
        in = 4'b1011; #20;
        in = 4'b1100; #20;
        in = 4'b1101; #20;
        in = 4'b1110; #20;
        in = 4'b1111; #20;

$display("Test Complete");
end
endmodule


